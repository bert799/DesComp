library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity memoriaROM is
   generic (
          dataWidth: natural := 13;
          addrWidth: natural := 9
    );
   port (
          Endereco : in std_logic_vector (addrWidth-1 DOWNTO 0);
          Dado : out std_logic_vector (dataWidth-1 DOWNTO 0)
    );
end entity;

architecture assincrona of memoriaROM is

  type blocoMemoria is array(0 TO 2**addrWidth - 1) of std_logic_vector(dataWidth-1 DOWNTO 0);

  function initMemory
        return blocoMemoria is variable tmp : blocoMemoria := (others => (others => '0'));
  begin
-- SETUP:
tmp(0):= "0100000000000000";	-- LDI R[0] $0
tmp(1):= "0101000000000000";	-- STA R[0] @0
tmp(2):= "0100010000000000";	-- LDI R[2] $0         	# Limpando o registrador das unidades
tmp(3):= "0100011000000000";	-- LDI R[3] $0         	# Limpando o registrador das dezenas
tmp(4):= "0100100000000000";	-- LDI R[4] $0         	# Limpando o registrador das centenas
tmp(5):= "0101000000001010";	-- STA R[0] @10        	# Espaço na memória dedicado ao milhar
tmp(6):= "0101000000001011";	-- STA R[0] @11        	# Espaço na memória dedicado à dezena de milhar
tmp(7):= "0101000000001100";	-- STA R[0] @12        	# Espaço na memória dedicado à centena de milhar
tmp(8):= "0100000000000001";	-- LDI R[0] $1
tmp(9):= "0101000000000001";	-- STA R[0] @1
tmp(10):= "0101000000000011";	-- STA R[0] @3         	# Utilizado para máscara de Bit menos significativo
tmp(11):= "0100000000001001";	-- LDI R[0] $9
tmp(12):= "0101000000000010";	-- STA R[0] @2         	# Comparação para definir o aumento do próximo HEX
tmp(13):= "0101000000010100";	-- STA R[0] @20        	# Redefinindo todos os HEX para 0
tmp(14):= "0101000000010101";	-- STA R[0] @21
tmp(15):= "0101000000010110";	-- STA R[0] @22
tmp(16):= "0101000000010111";	-- STA R[0] @23
tmp(17):= "0101000000011000";	-- STA R[0] @24
tmp(18):= "0101000000011001";	-- STA R[0] @25
tmp(19):= "0100000010000000";	-- LDI R[0] $128
tmp(20):= "0101000000000100";	-- STA R[0] @4         	# Utilizado para máscara de Bit mais significativo
tmp(21):= "0101000111111111";	-- STA R[0] @511       	# Limpando o botão de Incremento
tmp(22):= "0101000111111110";	-- STA R[0] @510       	# Limpando o botão de Alterar Limite
tmp(23):= "0101000111111011";	-- STA R[0] @507       	# Limpando o botão de RESET
tmp(24):= "0100000000000101";	-- LDI R[0] $5
tmp(25):= "0101000000000110";	-- STA R[0] @6         	# Comparção para minuto e segundo
tmp(26):= "0100000000000100";	-- LDI R[0] $4         	# Comparação para hora
tmp(27):= "0101000000000111";	-- STA R[0] @7
tmp(28):= "0100000000000010";	-- LDI R[0] $2
tmp(29):= "0101000000001000";	-- STA R[0] @8
-- # ========================================================= #
-- #                      LOOP PRINCIPAL                       #
-- # ========================================================= #
-- LOOP:
tmp(30):= "0001001101100000";	-- LDA R[1] @352
tmp(31):= "1011001000000011";	-- OPAND R[1] @3
tmp(32):= "1000001000000000";	-- CEQ R[1] @0         	# O botão de incremento não foi clicado
tmp(33):= "0111000000100100";	-- JEQ @TROCALIMITE
tmp(34):= "1001000000101010";	-- JSR @INCREMENTA
tmp(35):= "1001000001011011";	-- JSR @VERIFICA
-- TROCALIMITE:
tmp(36):= "0001001101100001";	-- LDA R[1] @353
tmp(37):= "1011001000000011";	-- OPAND R[1] @3
tmp(38):= "1000001000000000";	-- CEQ R[1] @0         	# O botão de troca de limite não foi clicado
tmp(39):= "0111000000011110";	-- JEQ @LOOP
tmp(40):= "1001000010010100";	-- JSR @SETLIMITE
tmp(41):= "0110000000011110";	-- JMP @LOOP
-- # ========================================================= #
-- #                     INCREMENTA VALOR                      #
-- # ========================================================= #
-- INCREMENTA:
tmp(42):= "0101000111111111";	-- STA @511
tmp(43):= "1000010000000010";	-- CEQ R[2] @2
tmp(44):= "1101000000000100";	-- RJEQ $4
tmp(45):= "0010010000000001";	-- SOMA R[2] @1
tmp(46):= "0101010100100000";	-- STA R[2] @288
tmp(47):= "1010000000000000";	-- RET         
tmp(48):= "0100010000000000";	-- LDI R[2] $0        	# Atualiza o dígito das dezenas
tmp(49):= "0101010100100000";	-- STA R[2] @288
tmp(50):= "1000011000000110";	-- CEQ R[3] @6
tmp(51):= "1101000000000100";	-- RJEQ $4
tmp(52):= "0010011000000001";	-- SOMA R[3] @1
tmp(53):= "0101011100100001";	-- STA R[3] @289
tmp(54):= "1010000000000000";	-- RET           
tmp(55):= "0100011000000000";	-- LDI R[3] $0        	# Atualiza o dígito das centenas
tmp(56):= "0101011100100001";	-- STA R[3] @289
tmp(57):= "1000100000000010";	-- CEQ R[4] @2
tmp(58):= "0111000000111110";	-- JEQ @ATMIL
tmp(59):= "0010100000000001";	-- SOMA R[4] @1
tmp(60):= "0101100100100010";	-- STA R[4] @290
tmp(61):= "1010000000000000";	-- RET
-- ATMIL:             	# Atualiza o dígito dos milhares
tmp(62):= "0100100000000000";	-- LDI R[4] $0
tmp(63):= "0101100100100010";	-- STA R[4] @290
tmp(64):= "0001101000001010";	-- LDA R[5] @10
tmp(65):= "1000101000000110";	-- CEQ R[5] @6
tmp(66):= "0111000001000111";	-- JEQ @ATDMIL
tmp(67):= "0010101000000001";	-- SOMA R[5] @1
tmp(68):= "0101101100100011";	-- STA R[5] @291
tmp(69):= "0101101000001010";	-- STA R[5] @10
tmp(70):= "1010000000000000";	-- RET
-- ATDMIL:            	# Atualiza o dígito das dezenas de milhar
tmp(71):= "0100101000000000";	-- LDI R[5] $0
tmp(72):= "0101101100100011";	-- STA R[5] @291
tmp(73):= "0101101000001010";	-- STA R[5] @10
tmp(74):= "0001101000001011";	-- LDA R[5] @11
tmp(75):= "1000101000000010";	-- CEQ R[5] @2
tmp(76):= "0111000001010001";	-- JEQ @ATCMIL
tmp(77):= "0010101000000001";	-- SOMA R[5] @1
tmp(78):= "0101101100100100";	-- STA R[5] @292
tmp(79):= "0101101000001011";	-- STA R[5] @11
tmp(80):= "1010000000000000";	-- RET
-- ATCMIL:            	# Atualiza o dígito das centenas de milhar
tmp(81):= "0100101000000000";	-- LDI R[5] $0
tmp(82):= "0101101100100100";	-- STA R[5] @292
tmp(83):= "0101101000001011";	-- STA R[5] @11
tmp(84):= "0001101000001100";	-- LDA R[5] @12
tmp(85):= "1000101000000010";	-- CEQ R[5] @2
tmp(86):= "0111000011011010";	-- JEQ @MAXOVERFLOW   	# Caso exceda o limite máximo do contador
tmp(87):= "0010101000000001";	-- SOMA R[5] @1
tmp(88):= "0101101100100101";	-- STA R[5] @293
tmp(89):= "0101101000001100";	-- STA R[5] @12
tmp(90):= "1010000000000000";	-- RET
-- # ========================================================= #
-- #                     VERIFICA LIMITE                       #
-- # ========================================================= #
-- ## A verificação começa com a centena de milhar
-- VERIFICA:
tmp(91):= "0001111000011001";	-- LDA R[7] @25
tmp(92):= "0011111000001100";	-- SUB R[7] @12
tmp(93):= "1011111000000100";	-- OPAND R[7] @4
tmp(94):= "1000111000000100";	-- CEQ R[7] @4
tmp(95):= "0111000011100111";	-- JEQ @OVERLIMIT
tmp(96):= "0001111000001100";	-- LDA R[7] @12
tmp(97):= "1000111000011001";	-- CEQ R[7] @25
tmp(98):= "0111000001100100";	-- JEQ @VERDMIL
tmp(99):= "1010000000000000";	-- RET
-- VERDMIL:
tmp(100):= "0001111000011000";	-- LDA R[7] @24
tmp(101):= "0011111000001011";	-- SUB R[7] @11
tmp(102):= "1011111000000100";	-- OPAND R[7] @4
tmp(103):= "1000111000000100";	-- CEQ R[7] @4
tmp(104):= "0111000011100111";	-- JEQ @OVERLIMIT
tmp(105):= "0001111000001011";	-- LDA R[7] @11
tmp(106):= "1000111000011000";	-- CEQ R[7] @24
tmp(107):= "0111000001101101";	-- JEQ @VERMIL
tmp(108):= "1010000000000000";	-- RET
-- VERMIL:
tmp(109):= "0001111000010111";	-- LDA R[7] @23
tmp(110):= "0011111000001010";	-- SUB R[7] @10
tmp(111):= "1011111000000100";	-- OPAND R[7] @4
tmp(112):= "1000111000000100";	-- CEQ R[7] @4
tmp(113):= "0111000011100111";	-- JEQ @OVERLIMIT
tmp(114):= "0001111000001010";	-- LDA R[7] @10
tmp(115):= "1000111000010111";	-- CEQ R[7] @23
tmp(116):= "0111000001110110";	-- JEQ @VERCEN
tmp(117):= "1010000000000000";	-- RET
-- VERCEN:
tmp(118):= "0101100000011110";	-- STA R[4] @30
tmp(119):= "0001111000010110";	-- LDA R[7] @22
tmp(120):= "0011111000011110";	-- SUB R[7] @30
tmp(121):= "1011111000000100";	-- OPAND R[7] @4
tmp(122):= "1000111000000100";	-- CEQ R[7] @4
tmp(123):= "0111000011100111";	-- JEQ @OVERLIMIT
tmp(124):= "1000100000010110";	-- CEQ R[4] @22
tmp(125):= "0111000001111111";	-- JEQ @VERDEZ
tmp(126):= "1010000000000000";	-- RET
-- VERDEZ:
tmp(127):= "0101011000011110";	-- STA R[3] @30
tmp(128):= "0001111000010101";	-- LDA R[7] @21
tmp(129):= "0011111000011110";	-- SUB R[7] @30
tmp(130):= "1011111000000100";	-- OPAND R[7] @4
tmp(131):= "1000111000000100";	-- CEQ R[7] @4
tmp(132):= "0111000011100111";	-- JEQ @OVERLIMIT
tmp(133):= "1000011000010101";	-- CEQ R[3] @21
tmp(134):= "0111000010001000";	-- JEQ @VERUNI
tmp(135):= "1010000000000000";	-- RET
-- VERUNI:
tmp(136):= "0101010000011110";	-- STA R[2] @30
tmp(137):= "0001111000010100";	-- LDA R[7] @20
tmp(138):= "0011111000011110";	-- SUB R[7] @30
tmp(139):= "1011111000000100";	-- OPAND R[7] @4
tmp(140):= "1000111000000100";	-- CEQ R[7] @4
tmp(141):= "0111000011100111";	-- JEQ @OVERLIMIT
tmp(142):= "1000010000010100";	-- CEQ R[2] @20
tmp(143):= "0111000010010001";	-- JEQ @LIMITE
tmp(144):= "1010000000000000";	-- RET
-- # =================== Chegou no limite ==================== #
-- LIMITE:
tmp(145):= "0100000011111111";	-- LDI R[0] $255
tmp(146):= "0101000100000000";	-- STA R[0] @256
tmp(147):= "0110000011101110";	-- JMP @END
-- # ========================================================= #
-- #                        SET LIMITE                         #
-- # ========================================================= #
-- SETLIMITE:
tmp(148):= "0101000111111110";	-- STA @510
tmp(149):= "0100000000000000";	-- LDI R[0] $0
tmp(150):= "0101000100100000";	-- STA R[0] @288
tmp(151):= "0101000100100001";	-- STA R[0] @289
tmp(152):= "0101000100100010";	-- STA R[0] @290
tmp(153):= "0101000100100011";	-- STA R[0] @291
tmp(154):= "0101000100100100";	-- STA R[0] @292
tmp(155):= "0101000100100101";	-- STA R[0] @293
tmp(156):= "0100110000000001";	-- LDI R[6] @1
tmp(157):= "0101110100000001";	-- STA R[6] @257
-- WAITUNI:
tmp(158):= "0001001101100001";	-- LDA R[1] @353
tmp(159):= "1011001000000011";	-- OPAND R[1] @3
tmp(160):= "1000001000000000";	-- CEQ R[1] @0
tmp(161):= "0111000010011110";	-- JEQ @WAITUNI
tmp(162):= "0101000111111110";	-- STA @510
tmp(163):= "0001110101000000";	-- LDA R[6] @320
tmp(164):= "0101110000010100";	-- STA R[6] @20
tmp(165):= "0101110100100000";	-- STA R[6] @288
-- WAITDEZ:
tmp(166):= "0001001101100001";	-- LDA R[1] @353
tmp(167):= "1011001000000011";	-- OPAND R[1] @3
tmp(168):= "1000001000000000";	-- CEQ R[1] @0
tmp(169):= "0111000010100110";	-- JEQ @WAITDEZ
tmp(170):= "0101000111111110";	-- STA @510
tmp(171):= "0001110101000000";	-- LDA R[6] @320
tmp(172):= "0101110000010101";	-- STA R[6] @21
tmp(173):= "0101110100100001";	-- STA R[6] @289
-- WAITCEN:
tmp(174):= "0001001101100001";	-- LDA R[1] @353
tmp(175):= "1011001000000011";	-- OPAND R[1] @3
tmp(176):= "1000001000000000";	-- CEQ R[1] @0
tmp(177):= "0111000010101110";	-- JEQ @WAITCEN
tmp(178):= "0101000111111110";	-- STA @510
tmp(179):= "0001110101000000";	-- LDA R[6] @320
tmp(180):= "0101110000010110";	-- STA R[6] @22
tmp(181):= "0101110100100010";	-- STA R[6] @290
-- WAITMIL:
tmp(182):= "0001001101100001";	-- LDA R[1] @353
tmp(183):= "1011001000000011";	-- OPAND R[1] @3
tmp(184):= "1000001000000000";	-- CEQ R[1] @0
tmp(185):= "0111000010110110";	-- JEQ @WAITMIL
tmp(186):= "0101000111111110";	-- STA @510
tmp(187):= "0001110101000000";	-- LDA R[6] @320
tmp(188):= "0101110000010111";	-- STA R[6] @23
tmp(189):= "0101110100100011";	-- STA R[6] @291
-- WAITDMIL:
tmp(190):= "0001001101100001";	-- LDA R[1] @353
tmp(191):= "1011001000000011";	-- OPAND R[1] @3
tmp(192):= "1000001000000000";	-- CEQ R[1] @0
tmp(193):= "0111000010111110";	-- JEQ @WAITDMIL
tmp(194):= "0101000111111110";	-- STA @510
tmp(195):= "0001110101000000";	-- LDA R[6] @320
tmp(196):= "0101110000011000";	-- STA R[6] @24
tmp(197):= "0101110100100100";	-- STA R[6] @292
-- WAITCMIL:
tmp(198):= "0001001101100001";	-- LDA R[1] @353
tmp(199):= "1011001000000011";	-- OPAND R[1] @3
tmp(200):= "1000001000000000";	-- CEQ R[1] @0
tmp(201):= "0111000011000110";	-- JEQ @WAITCMIL
tmp(202):= "0101000111111110";	-- STA @510
tmp(203):= "0001110101000000";	-- LDA R[6] @320
tmp(204):= "0101110000011001";	-- STA R[6] @25
tmp(205):= "0101110100100101";	-- STA R[6] @293
-- # ============ Retornando o valor do contador ============= #
tmp(206):= "0101010100100000";	-- STA R[2] @288
tmp(207):= "0101011100100001";	-- STA R[3] @289
tmp(208):= "0101100100100010";	-- STA R[4] @290
tmp(209):= "0001101000001010";	-- LDA R[5] @10
tmp(210):= "0101101100100011";	-- STA R[5] @291
tmp(211):= "0001101000001011";	-- LDA R[5] @11
tmp(212):= "0101101100100100";	-- STA R[5] @292
tmp(213):= "0001101000001100";	-- LDA R[5] @12
tmp(214):= "0101101100100101";	-- STA R[5] @293
tmp(215):= "0100110000000000";	-- LDI R[6] @0
tmp(216):= "0101110100000001";	-- STA R[6] @257
tmp(217):= "1010000000000000";	-- RET
-- # ========================================================= #
-- #                         OVERFLOW                          #
-- # ========================================================= #
-- MAXOVERFLOW:
tmp(218):= "0100010000001001";	-- LDI R[2] $9
tmp(219):= "0100011000001001";	-- LDI R[3] $9
tmp(220):= "0100100000001001";	-- LDI R[4] $9
tmp(221):= "0101010000001010";	-- STA R[2] @10
tmp(222):= "0101010000001011";	-- STA R[2] @11
tmp(223):= "0101010000001100";	-- STA R[2] @12
tmp(224):= "0101010100100000";	-- STA R[2] @288
tmp(225):= "0101010100100001";	-- STA R[2] @289
tmp(226):= "0101010100100010";	-- STA R[2] @290
tmp(227):= "0101010100100011";	-- STA R[2] @291
tmp(228):= "0101010100100100";	-- STA R[2] @292
tmp(229):= "0101010100100101";	-- STA R[2] @293
tmp(230):= "0110000011101010";	-- JMP @OVERFLOW
-- OVERLIMIT:
tmp(231):= "0100000011111111";	-- LDI R[0] $255
tmp(232):= "0101000100000000";	-- STA R[0] @256
tmp(233):= "0110000011101010";	-- JMP @OVERFLOW
-- OVERFLOW:
tmp(234):= "0101000111111111";	-- STA @511
tmp(235):= "0100000000000001";	-- LDI R[0] $1
tmp(236):= "0101000100000010";	-- STA R[0] @258
tmp(237):= "0110000011101110";	-- JMP @END
-- # ========================================================= #
-- #                         LOOP END                          #
-- # ========================================================= #
-- END:
tmp(238):= "0001001101100100";	-- LDA R[1] @356
tmp(239):= "1011001000000011";	-- OPAND R[1] @3
tmp(240):= "1000001000000001";	-- CEQ R[1] @1
tmp(241):= "0111000011110111";	-- JEQ @CLEAR
tmp(242):= "0001001101100000";	-- LDA R[1] @352
tmp(243):= "1011001000000011";	-- OPAND R[1] @3
tmp(244):= "1000001000000001";	-- CEQ R[1] @1
tmp(245):= "0111000011101010";	-- JEQ @OVERFLOW
tmp(246):= "0110000011101110";	-- JMP @END
-- # ========================================================= #
-- #                          CLEAR                            #
-- # ========================================================= #
-- CLEAR:
tmp(247):= "0100000000000000";	-- LDI R[0] $0
tmp(248):= "0101000100100000";	-- STA R[0] @288
tmp(249):= "0101000100100001";	-- STA R[0] @289
tmp(250):= "0101000100100010";	-- STA R[0] @290
tmp(251):= "0101000100100011";	-- STA R[0] @291
tmp(252):= "0101000100100100";	-- STA R[0] @292
tmp(253):= "0101000100100101";	-- STA R[0] @293
tmp(254):= "0101000100000000";	-- STA R[0] @256
tmp(255):= "0101000100000001";	-- STA R[0] @257
tmp(256):= "0101000100000010";	-- STA R[0] @258
tmp(257):= "0101000111111111";	-- STA R[0] @511
tmp(258):= "0101000111111110";	-- STA R[0] @510
tmp(259):= "0101000111111011";	-- STA R[0] @507
tmp(260):= "0110000000000000";	-- JMP @SETUP




		return tmp;
    end initMemory;

    signal memROM : blocoMemoria := initMemory;

begin
    Dado <= memROM (to_integer(unsigned(Endereco)));
end architecture;